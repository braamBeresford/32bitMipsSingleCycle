module topLevel ();


endmodule