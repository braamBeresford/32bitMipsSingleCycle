module topLevel();


endmodule