module topLevel ();


endmodule