module topLevel();



end module